module bondpad_70x70_novias (
    inout pad
);
endmodule
